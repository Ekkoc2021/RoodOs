� ��  � ��� �   �� tO�� tJ�ú�����B� B�B��B� B�f1ۈ�f�   � ������$�<u󐐐���&�GG��K�� u��                                                                                                                                                                                                                                                                                                                                                                                                                 U��T'  �'           ��   �� ��   ��                                                 f1�f�PAMS��f� �  f�   �χ���f�� u���� �f��"�f�   f� �؎��Ў�༠  �  ���
   �   �    �   � 0  �u   � 0  ��� ,  �    �   � 0  �    �   ����	���   ���E ���  �� �� ��    "� �   �"� � ���"�� � Q�   � ��Y�f������fB�f����fB�f����fB�f����$�fB� fB�1ۈ˹   f� ���f���$�<u򐐐f��f�&f�GG��K�� u��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       f� �؎��Ў�� � ��    �   �R�    P�   �PQS��0  ��PR1�1�f����f����f����f����ZX�RPf����f�����f����f�����XZ�U����]�U����Ef�E��E�U�P�E�U�f��E�U�P���U����Ef�E�E�E��E�E�f�E�  �"�U��E���M��U��� ��E���f�E��E�f;E�rԐ���U����E�@9Er�    �>�E� ���U�E��E�@�E��E� ���M��U��P�uR�a������   ��U����E�@9Er�    �-�E� ���U�E��E�@�E��U��E�E��   ��U����E�@��u�E�@���u�E�@�E�E�E��E�    �E�   �H�E� ���E�E�Ѓ��u�P�E�Ѓ���~�E� ���E�E�ЉE�E�E��E��E�@9E�r��E���U��E�U��E��    �E�P�E�@    �]�U��E�U��E�U�P�E�@    �]�U����E� �E��E���   ����ЈE��E���E�E��E��� �U�
�U��
E���E�@�P�E�P��U����E� �E��E���   ������ЈE��E���E�E��E��� �U�
�U��"E���E�@�P��E�P��U��� �E�@    �E� �E�E�@���E��E�    ��E���    �E���     �E��E�@���E�9�wՋE�@���E��E�    � �E��E���    �E�ȃ���  �E��E���9E�|Ր���U��S���E�@9Er�   �=�E��E���� �E��U��E���   �����!E�������ЈE��E��]���U��� �E� �E�E�@�����E��E�    �%�E���    �E�Ћ ���t�E����E���E��E�@���E�9�w��E�    �E�@����u�E�@���E���E�@�����E�E��E��z�E��E��� <�te�E�    �V�E���    �E��P�u���������u3�E���    �E�ЉE�@9�r������0�E���    �E����E��}�~��E��E�9E��z����������U��� �E� �E��E�@�����E��E�    �E�@����u�E�@�����E���E�@���E��E��E��v�E��E��� <�ta�E�   �R�E��    �E�ЉE�@9�s3�E��    �E��P�u���������u�E��    �E����   �m��}� y��m��E��P��E�9��y����E�    �%�E��    �E�Ћ ���t�E����E���E��E�@���E�9�wɋE�@�����E��s�E��E��� <�t^�E�   �O�E��    �E�ЉE�@9�s0�E��    �E��P�u��������u�E��    �E��� �m��}� y��m��E��P��E�9�r��������U��� �E� �E�E�@�����E��E�    �$�E���    �E�Ћ ��t�E����E���E��E�@���E�9�w��E�    �E�@����u�E�@���E���E�@�����E�E��E��s�E��E��� ��t^�E�    �O�E���    �E��P�u��������t,�E���    �E�ЉE�@9�s�E���    �E����E��}�~��E��E�9E�w��������U��� �E� �E��E�@�����E��E�    �E�@����u�E�@�����E���E�@���E��E��E��v�E��E��� ��ta�E�   �R�E��    �E�ЉE�@9�s3�E��    �E��P�u��������t�E��    �E����   �m��}� y��m��E��P��E�9��y����E�    �$�E��    �E�Ћ ��t�E����E���E��E�@���E�9�wʋE�@�����E��s�E��E��� ��t^�E�   �O�E��    �E�ЉE�@9�s0�E��    �E��P�u�<�������t�E��    �E��� �m��}� y��m��E��P��E�9�r��������U���   �E� P��E�    �0�E���E��� ��t����U�ʈ�E���E�E��}�w�} u����}� u�E� 0�E���  �;�U�E���  �E�    ��E�+E����M�U����t�����E��E�;E�r���U���   �E� P��E��E�    �0�E���E��� ��s����U�ʈ�E���E�E��}�w�} u����}� y
�E� -�E�}� u�E� 0�E���  �;�U�E���  �E�    ��E�+E����M�U����s�����E��E�;E�r���U����E�    ��U�E�ЋM�U��� ��E��E�;Erߐ���U����E�E��E�    �U�E��� ��u�������U�E��� 8E�u�E���E�����U����E�    �U�E����M�E��� 8�t �U�E��� ���U�E��� ��)���U�E��� ��u�    ��E����U����E�    ��E��U�E��� ��u�E���U����E�    ��U�E�ЋM�U��� ��E��E�;ErߋU�E���  �E��U����E�    ��U�E�ЋM�U��� ��E��U�E��� ��u؋U�E���  �E���U����u�D������E��E�    ��U�E�ЋM�U��� ��E��E��E�;ErۋU�E���  �E��U���8�E� �E�    �U�E��� < t%�U�E��� <-u�u���U�E��� <+u��E��Ɛ�E�E�E�    ���]���E��XP����]�E��U�E��� ��t�U�E��� </~�U�E��� <9~����]��E�    �4�E��XP����]�U�E��� ����0�E��E��M��E����]��E��E�;E�rċU�E��� <.t�}� t
�E����   �E��   �E��E�E�    �4�E��XP����]�U�E��� ����0�E��E��M��E����]��E��U�E��� ��t�U�E��� </~�U�E��� <9~��}� t�E�����E���U��� �E� �E�    �U�E��� < t%�U�E��� <-u�u���U�E��� <+u��E��Ɛ�E�E�E�    �E�   ��U��������E��E��U�E��� ��t�U�E��� </~�U�E��� <9~��E�    �E�    �.�E�����������E��U�E��� ����0�E�E�E��E�;E�rʀ}� t�E�����E���U���8�E�E��E�E��E��}��Eހ�f�E��m��}��mދEЉE�E��    �EЉU��m��E����]��E��P�u�  ���E�U�E��� .�E�    �E�������v�E����]��E�   �}��Eހ�f�E܃E��E��XP����]��E��m��}��mދEЉE�E�H0�U�E�Љʈ�E�    �EЉU��m��E����]��} t�E�;Es+�} u�E�������z�E�������t�}�w
�E��x�����E�P�E��  �E���U����E� �E�   �E�E���E��E������������E��}� u�}� t
�E� -�E�U�E���  �E�    �G�M����̉�����������)��ʉЍP0�E�+E�H��EȈ�E�����������E�E��E�;E�r��}� t�E�����E���U��S���E� �} y�E��]�E�   �E�E���E��E�����������E��}� u�}� t
�E� -�E�U�E���  �E�    �[�M�gfff�����������)؉�����)��ʉЍP0�E�+E�H��EȈ�M�gfff�����������)ЉE�E��E�;E�r��}� t�E����E�]���U���h�E�E��E�    �E�    �  �U�E�� <%t�U�EЋM��U�� ��b  �E�P�E�� �E��E��c���+  ��P����E��E܍P�U܋ P�E�P�������U��EE�PR�g������U�Ѓ��E���   �E��E܍P�U�� �]�j �u��u��E�P�Y������U��E��E�PR�������U�Ѓ��E��   �E��E܍P�U܋ �M��Uʃ�PR��������U�Ѓ��E��x�E��E܍P�U܋�M��EȈ�]�E��E܍P�U܋P� ��P�E�P��������U��E��E�PR�������U�Ѓ��E���U�EЋM��U�� ���E��E��U�E�� ���Z����U��E��  �E���U����E�E��E�    ��U�E���E��E��E�;Er搐��U�����h`P��l  �����uhvP��Y  �����uh�P��F  �����uh�P��3  �����uh�P��   ��������U�����h�P��  �����U�����h�P���  �����U��S���E�X�E�H�E��E�@��SQRPh�P��  �� ��]���U��S��   �E� � ����PhQ��  ��f�E�  �
  �E� �H�U��������ȋ ����p���RP��������E� �H�U��������ȋ ��P��p���Ph1Q��  ���E� �H�U��������ȋ@��PhBQ���  ���E� �H�U��������ȋ@��PhWQ���  ���E� �H�U��������ȋP�E� �X�M��������؋@��RPhhQ��  ���E���f�E��E� � f9E�������E�H�E�P�E�@��QRPh�Q��<  ���E�    �Q�E�P���u���l���PR�������E�P�E���Ѓ�Ph�Q���  ����l�����P�������E��E�@9E�r����]���U��VS���   ��h�Q��  ����d� 0��E�H�E��������ȣ�d���d�f�   ��d���d����P�E�    �E� ��PhR��W  ��f�E�  �E�    f�E�  �I  �E�H�U�������ȋP� ����Z���PR�������E�H�U�������ȋP� RP��Z���Ph1Q���  ���E�H�U�������ȋP�@��RPhR��  ���E�H�U�������ȋ@��Ph)R��  ���E�H�U�������ȋ@���c  �E�H�U�������ȋP� f%�f�E�f�}� ��   �E�H�U�������ȋP�    �� ���ӋE�p�U�������Ɖȉ�������V�E�H�U�������ȋH�X�Uڸ   )Љ�@���������D����E�p�U�������Ɖȉ�+�@����D����F�V��d����f��E�H�U�������ȋ�X��d��p��d�� �Љ����������ʉ�E�H�U�������ȋP�@�á�d��H��d�� �Љ��������ȁ� ����ډP��d��H��d�� �Љ��������ȋH��d��X��d�� �Љ������������ʉP��d��H��d�� �Љ����������E��B��d��H��d�� �Љ��������ȋ@E��d��H��d�� �Љ��������ȋU����P�E�H�U�������ȋP�@E��E��f�E��U�E� 9���������u��u�h8R���  ���E��d���d�    f��d� �E�����u�E����	�E������E���d��E�ЉE܋Eܣ�d���d�    �E�    �`��d��E���
Ѓ�Ph    ��H�����P�������E�����H�����d�����d����u荅H���Ph�d��%������E��E���
9E�r��E�%�  ��tm��d�����H�����d���d���
E�%�  ����RP��H�����P�#�������d�����d���d�����P��H���Ph�d���������htR��y  ����d��e�[^]�U���(�E�H�E�P�������ȉE��E�%�  ��u�E�   @����E�   @�����E���u�h�R��  ���E�   @��P�u�  ���E�E� �H�U�������ȋ ��P�u��   ���E�E�P���u�E�PR�������E�    �(�E������u�P�!������E�@�P�E�P�E��E�;E�rЋE�����U��S���E�E��E�E�E��P�E��@��)��E�P�E�X��)�9�v�   �0�E��P�E��@��)��E�P�E�X��)�9�s�������    �]���U����E� �@�E��E�    �A�U���������E�Ћ@9Er!�U���������E�Ћ@9Ew�E���E��E� � ��9E�r��E� � ����U��S��$�E���E��h|-��u��������E��E�@9E�rh�R�h�R�h�   h�R����������u��E�P�u��������E��P�E��@9�u
�    �   �E����E���u��)������E�� ЉE���u��u��c������E�@�P�E�P���u��u�������E�E� �H�U�������ȋ�E� �X�U�������؋P�E�)���ȋ]���U����E� �@�E��E�    �X�U���������E�Ћ 9Er9�U���������E�Ћ�U���������E�Ћ@�9Es�E���E��E� � ��9E�r��E� � ����U��S��$�E% ����E��u��u�T������E��E� �H�U��������ȋ�E�)����ËE� �H�U��������ȋ@؉E�E����E�E�P�E���Ѓ��E�E� �H�U��������ȋP�E�)Ѓ�P�u��������E�@�P��E�P��]���U��S��$f�E�  �  �E��U�R�� ��PR�����������   �E�f ����P�u�$  ��% ����E��E�f ����P�u��  �����E�f ����P�u��  ���U�SPRh�R��|  ��f�E� �E�    �_�E�����P�u��  ���E܃}� t=�E��f�E���u��u�hS��.  ���E��f��u��h(S��  ���E��}��  v��E���f�E�f�}�� �����f�E�  ��   �E��P�u�&  ��% ����E��E�U�R��`��PR����������   �E��P�u��   �����E��P�u��  ���U�SPRh�R��j  ��f�E� �E�    �b�E������P�u��  ���E��}� t=�E��f�E���u��u�h*S��  ���E��f��u��h(S���  ���E��}��  v��E��f�E�f�}���������]���U����Ef�E�E�@��,�E�f�}��v�E� ��� �E��� ����E�@��l�E��E� �E��� ����U���(�Ef�E��E��P�u�  ��% ����E��Ef�E�� �E���Pj �u��$  ���E���f�E�f�}�� v�f�E�  � �E��j�P�u�  ���E��f�E�f�}��v؋E�����E��RP�u��  ���i   �E�-   �E�@�� ��RP�;��������U��E8�]�U����E% ������E��E� 0 ��E����  �E��h �?�����������U����E� 0 ��E��  � ��  ���U����u�������E� �?���h   j �u��h������������U����Ef�E��u�_������E� �?��E��    �E�E��t������U���(�Ef�E�E�@�E��E��    �E�E�f�}��v#�E�-   �E�@�� ��RP��������E�U�R��`��PR���������U���(�Ef�E�E�@�E��E��    �E���     f�}��v=�E�-   �E�@�� ��RP��������E�@�U��   ��f�DP���.�E�U�R��`��PR�������E�@�U��0f�DP����U����Ef�E��u�������E� �?��E��    �E�Ћ �E��%����E���U����U�Ef�U�f�E�f�}��v;�E�@�U���   ���DP���E���E�@�U���   ��f�LP�-�E�@�U���0�DP���E���E�@�U���0f�LP��U����U�Ef�U�f�E�f�}��v�E�@�U���   �J�U�f�TH��E�@�U��J0�U�f�TH��U����Ef�E�E�@�E��E��    �E�Ћ ��U����u��������E� �?�f�E�  �(�E���    �E�Ћ 9Eu�E���E���f�E�f�}��v�������   ��U����E�e��E� e��e� e��E�e��e��¡e��� ��Rh   P�K������e��¡e���`��Rh   P�*������ e���U����E�@�� ��P�������f ��U���f�E�  �D�E�@�U����DPf��x"�E�@�U����DPf=�
�E�f ��E���f�E�f�}�� v��   ��U���:�E�@�Lg��҃��DPf��u�Lg�f �8�Lg���f�Lg��Lg�f=� ~��Lg�f= u	f�Lg�  �   ]�U����E�@��`��P���������U���f�E�  �@�E�@�U���0�DPf��x�E�@�U���0�DPf=��E���E���f�E�f�}��v��   ��U���6�E�@�Ng��҃�0�DPf��u	�Ng��8�Ng���f�Ng��Ng�f=�~��Ng�f= u	f�Ng�  �   ]�U���   �E�pg��E�lg���h8S���  �����uh\S��  ���U�EЃ�Ph�S��  ����hlg��������E�U�EЃ�h�g��uP�D������E��hg��7��E��`g��E�dg����u����������u���������E�E�    ��P�����T���߭P�����S������d$��$h�S���  �����u��9�����f�E� �E��Ph�S���  ���E�U�����PR�u��:��������u���������h�S��  ����h`g��)   ���E���u�����������u��J������`g���U���(�8����E� ��P�������E��}� u
�    �  �E�@��P�p�����f�E�f�}� ��   �E�@��P�1�����f�E�f�}��u�E� ���u�P��������    �E  �E� ��P�=������E�}� u�E� ���u�P��������    �  ���u��F������E��ЋE�����E�@��RQP�������E��ЋE�@��j RP�O������E��ЋE�@��RP������% ����E��j �u�������f�E�f�}��v�E� ���u�P�������    �g�E�U�����PR�u���������E��ЋE�@��jRP�:����������E������E���ЉE��E���P������������E���U���(�e����E� ��P��������E��}� u
�    �  �E�@��P������f�E�f�}� ��   �E�@��P�s�����f�E�f�}��u�E� ���u�P�)������    �@  �E� ��P�j������E�}� u�E� ���u�P��������    �  ���u��s������E��ЋE�����E�@��RQP��������E��ЋE�@��j RP�|������E��ЋE�@��RP������% ����E��j �u��������f�E�f�}��v�E� ���u�P�H������    �b�E�U�����PR�u���������E��ЋE�@��jRP�g������E������E���ЉE��E���P������������E���U��������E���E�E��%�  �E��E��ЋE�@��RP����������E�E�����P�u����������E�E� ���u�P�m������E����U�R��Pj R�!������E��ЋE�@��j�RP�������������U����c�U��E�@��RP�D�����% ����E��E� ���u�P��������U��E�@��j�RP�������U��E�@��RP�A������E�@��P�_�����f�E�f�}���{����c�U��E�@��RP������% ����E��E� ���u�P�m������U��E�@��j�RP�6������U��E�@��RP�������E�@��P������f�E�f�}���{������ÍL$����q�U��VSQ���ˋC� ���Ph�S���   ���C��� ��Ph	T��   ���'   �s�K�S�VQRP�������    �e�Y[^]�a��U��S����h T��l   ����m�@T���m�GT���m�  ��m� ���hMT��4   ����m���m���m���m���SQRPhdT��	   �� ��]���U���h�E�E��E�    �Q  �U�E�� <%t�U�E�� ����P��  ���  �E�P�E�� �E��E��c����   ���T����E��E�P�U� ��P�E�P���������E�P�v  ����   �E��E�P�U�� �]�j �u��u�E�P����������E�P�<  ���   �E��E�P�U� ��P�������k�E��E�P�U� ����P�  ���K�E��E�P�U� ���U�RP���������E�P��  ����U�E�� ����P��   ����E��U�E�� �����������U����} u�E��0��P�   ���   �E� �E� ʚ;�E� �E�    �c�E��}��E�E��}��U�}� u
�}� t�E��}� t�E��0�E��E��P�*   ���M�gfff�����������)ЉE��E��}�	~���U���(�E�E��E�E��E� ���E�P��   �����U�����  �E�M��gfff�����������)ЉE��E�    ��"   �m�P���u���  ���E��E�;E�|ݐ���U����E� ��f�E�� f�E�  �  ��E��E�    �1�U��E���M�U��� ��E���f�E��E��f�E�E��E�;E�|ǐ���U����E� ���E�    �  ��E��E�    �U�E�� ����   �U�E�� <uF�M�gfff���������)ȉ�������E��E����������P��   ���E��   �U�E�� <
u[�M�gfff�����������)ЉE�}�u	������m��E�P��������E��E����������P�g   ���E��5�U�EЋM��U��� ��E��E����������P�0   ���E����������U��S���E�    ������؉E�E�]���U��S���E���������]���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          0123456789ABCDEF    �#��"��#�#��#��#��#��#��#��#��#��#��#��#��#��#�c#�      $@


!!!!! error !!!!!
 filename:%s 
 line:%d 
 function:%s 
 condition:%s 
 disallowInterrupt!!!!!!
 enableInterrupt!!!!!!
    indexBitsAddr:0x%p,indexOfBitMap:%d,size:%d,used:%d
 Block of available memory:%d
   addr: 0x%s\%d    memory size: %d B    bitsize: %d 
       bitIndex between %d and %d 
   indexLisnt:elementSize: %d length :%d dataAddr: 0x%p 
    data details  addr:0x%p
      Physical memory initialization...
 Block of memory:%d
   size: %d B    type: %d 
     total available memory : %d Byte ,total bitmap size : %d
 Physical memory Initialization successful!
 size of the kernel: %d Page 
 index < list->length  src/kernel/memory/physicalMem.c getPhyPage index:%d,PDE:0x%p,PTSzie:%d 
  %d :0x%p  
  %d :%p       Init memory management module...
   pageTable physical addr : 0x%p 
    pageTable virtual addr : 0x%p 
 The kernel uses memory size: %f KB! 
   the index of kernel pde : %d 
 
              �@gdt   count:%d 
 gdt virtual addr:0x%p
 Kernel was loaded successful !
 RoodOs 0.0.1 Welcom to RoodOs! ^_^
 ___%s__%s_ 
kernel p\v addr:0x%p\0x%p
  �B�YB�3C��B�3C�3C�3C�3C�3C�3C�3C�3C�3C�C�3C�3C��B�